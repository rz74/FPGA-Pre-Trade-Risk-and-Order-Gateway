`timescale 1ns/1ps
// Apply post-decision state changes (positions, credit usage, CAM/STP entries).
module state_update (
    input  wire clk,
    input  wire rst_n
    // TODO: inputs: decision + order fields; side-effects into BRAM/CAM
);
// TODO
endmodule
