`timescale 1ns/1ps
// AXI-Lite register block for config plane (limits, collars, kill-switch, status).
module axi_lite_regs (
    input  wire clk,
    input  wire rst_n
    // TODO: AXI-Lite interface; register map TBD
);
// TODO
endmodule
