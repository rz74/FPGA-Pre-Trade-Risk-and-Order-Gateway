`timescale 1ns/1ps
module snapshot_mux (
    input  wire clk,
    input  wire rst_n
    // TODO: route NBBO/limits snapshots to checks (per-symbol/account)
);
// TODO
endmodule
