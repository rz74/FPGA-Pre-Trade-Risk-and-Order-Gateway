`timescale 1ns/1ps
// Check #3/4: credit/exposure and position limits
module credit_position_check (
    input  wire clk,
    input  wire rst_n
    // TODO: inputs: account, symbol, qty, notional; outputs: pass/fail + reason
);
// TODO
endmodule
