`timescale 1ns/1ps
// Simple per-symbol NBBO cache (bid/ask/ts). Backed by BRAM.
module nbbo_cache (
    input  wire clk,
    input  wire rst_n
    // TODO: write port for ITCH-derived updates; read port for checks
);
// TODO
endmodule
