`timescale 1ns/1ps
// Check #1: max order size & notional
module size_notional_check (
    input  wire clk,
    input  wire rst_n
    // TODO: inputs: qty, price (from order + NBBO); outputs: pass/fail + reason code
);
// TODO
endmodule
