`timescale 1ns/1ps
module account_limits_bram (
    input  wire clk,
    input  wire rst_n
    // TODO: credit/exposure, per-account limits; atomic updates
);
// TODO
endmodule
