`timescale 1ns/1ps
module ingress_unpack (
    input  wire clk,
    input  wire rst_n
    // TODO: s_axis_order_intent, field extraction
);
// TODO
endmodule
