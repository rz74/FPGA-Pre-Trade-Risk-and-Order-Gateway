`timescale 1ns/1ps
// Check #2: price collar vs NBBO
module price_collar_check (
    input  wire clk,
    input  wire rst_n
    // TODO: inputs: order side/price, NBBO; configurable collar bps
);
// TODO
endmodule
