`timescale 1ns/1ps
// Check #5: token-bucket throttling (message-rate cap)
module throttle_bucket (
    input  wire clk,
    input  wire rst_n
    // TODO: parameters: refill rate, burst; input: order pulse; output: allow/drop
);
// TODO
endmodule
