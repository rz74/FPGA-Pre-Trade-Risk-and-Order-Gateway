`timescale 1ns/1ps
// Check #6: duplicate order ID prevention via small CAM
module dupid_cam (
    input  wire clk,
    input  wire rst_n
    // TODO: lookup+insert order_id; eviction by epoch
);
// TODO
endmodule
