`timescale 1ns/1ps
module symbol_limits_bram (
    input  wire clk,
    input  wire rst_n
    // TODO: per-symbol max size, price collar %, position caps
);
// TODO
endmodule
