`timescale 1ns/1ps
// Epoch counter/ticker for time-based eviction in CAM/STP/throttle
module epoch_ctrl (
    input  wire clk,
    input  wire rst_n
    // TODO: parameters: tick period; outputs: epoch number
);
// TODO
endmodule
